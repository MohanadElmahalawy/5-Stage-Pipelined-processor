library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
ENTITY CCR IS
PORT
(
	CLK:IN STD_LOGIC;
	FLAGS_IN :IN STD_LOGIC_VECTOR(2 DOWNTO 0); --- Z N C---
	Enablee: IN STD_LOGIC;
	FLAGS_OUT:OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
	RESET_Z:IN STD_LOGIC;
	RESET_N:IN STD_LOGIC;
	RESET_C:IN STD_LOGIC;
	RESET:IN STD_LOGIC;
	SET_C:IN STD_LOGIC;
	SET_CCR:IN STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END ENTITY CCR;
ARCHITECTURE CCR_ARCH OF CCR IS 
	SIGNAL TEMP_FLAG : STD_LOGIC_VECTOR(2 DOWNTO 0);
BEGIN
	PROCESS (CLK, Enablee,RESET_Z,RESET_N,RESET_C,SET_C,RESET)
	BEGIN
		IF RESET_Z='1' THEN
			TEMP_FLAG(2)<='0';
		ELSIF RESET_N='1' THEN
			TEMP_FLAG(1)<='0';
		ELSIF RESET_C='1' THEN
			TEMP_FLAG(0)<='0';
		ELSIF RESET='1' THEN
			TEMP_FLAG<="000";
		ELSIF RISING_EDGE(CLK)  THEN
			IF Enablee='1' THEN
				IF SET_C='1' THEN
					TEMP_FLAG(0)<='1';
				ELSE 
					TEMP_FLAG<=SET_CCR;
				END IF;
			ELSE 
				TEMP_FLAG<=FLAGS_IN;
			END IF;
		END IF;
	END PROCESS;
	FLAGS_OUT<=TEMP_FLAG;
END CCR_ARCH;